Miraculous Treasure
ds
